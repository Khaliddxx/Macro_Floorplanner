#N
addr[0], LAYER met3 ( -2000 -300 ) ( 2000 300 )
addr[1], LAYER met3 ( -2000 -300 ) ( 2000 300 )
addr[2], LAYER met2 ( -140 -2000 ) ( 140 2000 )
addr[3], LAYER met2 ( -140 -2000 ) ( 140 2000 )
addr[4], LAYER met2 ( -140 -2000 ) ( 140 2000 )
addr[5], LAYER met2 ( -140 -2000 ) ( 140 2000 )
addr[6], LAYER met3 ( -2000 -300 ) ( 2000 300 )
config_in[0], LAYER met2 ( -140 -2000 ) ( 140 2000 )
config_in[1], LAYER met2 ( -140 -2000 ) ( 140 2000 )
config_in[2], LAYER met3 ( -2000 -300 ) ( 2000 300 )
config_in[3], LAYER met2 ( -140 -2000 ) ( 140 2000 )
config_in[4], LAYER met2 ( -140 -2000 ) ( 140 2000 )
config_in[5], LAYER met2 ( -140 -2000 ) ( 140 2000 )
config_in[6], LAYER met2 ( -140 -2000 ) ( 140 2000 )
config_in[7], LAYER met2 ( -140 -2000 ) ( 140 2000 )
#S
config_out[0], LAYER met2 ( -140 -2000 ) ( 140 2000 )
config_out[1], LAYER met3 ( -2000 -300 ) ( 2000 300 )
config_out[2], LAYER met3 ( -2000 -300 ) ( 2000 300 )
config_out[3], LAYER met3 ( -2000 -300 ) ( 2000 300 )
config_out[4], LAYER met2 ( -140 -2000 ) ( 140 2000 )
config_out[5], LAYER met2 ( -140 -2000 ) ( 140 2000 )
config_out[6], LAYER met3 ( -2000 -300 ) ( 2000 300 )
config_out[7], LAYER met2 ( -140 -2000 ) ( 140 2000 )
out, LAYER met3 ( -2000 -300 ) ( 2000 300 )
#E
config_clk, LAYER met3 ( -2000 -300 ) ( 2000 300 )
config_en, LAYER met2 ( -140 -2000 ) ( 140 2000 )