#N
x[0], LAYER met3 ( -2000 -300 ) ( 2000 300 )
x[1], LAYER met3 ( -2000 -300 ) ( 2000 300 )
x[2], LAYER met3 ( -2000 -300 ) ( 2000 300 )
x[3], LAYER met3 ( -2000 -300 ) ( 2000 300 )
x[4], LAYER met3 ( -2000 -300 ) ( 2000 300 )
x[5], LAYER met2 ( -140 -2000 ) ( 140 2000 )
x[6], LAYER met2 ( -140 -2000 ) ( 140 2000 )
x[7], LAYER met2 ( -140 -2000 ) ( 140 2000 )
x[8], LAYER met3 ( -2000 -300 ) ( 2000 300 )
x[9], LAYER met2 ( -140 -2000 ) ( 140 2000 )
x[10], LAYER met2 ( -140 -2000 ) ( 140 2000 )
x[11], LAYER met2 ( -140 -2000 ) ( 140 2000 )
x[12], LAYER met3 ( -2000 -300 ) ( 2000 300 )
x[13], LAYER met3 ( -2000 -300 ) ( 2000 300 )
x[14], LAYER met3 ( -2000 -300 ) ( 2000 300 )
x[15], LAYER met2 ( -140 -2000 ) ( 140 2000 )
x[16], LAYER met2 ( -140 -2000 ) ( 140 2000 )
x[17], LAYER met2 ( -140 -2000 ) ( 140 2000 )
x[18], LAYER met2 ( -140 -2000 ) ( 140 2000 )
x[19], LAYER met3 ( -2000 -300 ) ( 2000 300 )
x[20], LAYER met2 ( -140 -2000 ) ( 140 2000 )
x[21], LAYER met3 ( -2000 -300 ) ( 2000 300 )
x[22], LAYER met2 ( -140 -2000 ) ( 140 2000 )
x[23], LAYER met3 ( -2000 -300 ) ( 2000 300 )
x[24], LAYER met2 ( -140 -2000 ) ( 140 2000 )
x[25], LAYER met2 ( -140 -2000 ) ( 140 2000 )
x[26], LAYER met2 ( -140 -2000 ) ( 140 2000 )
x[27], LAYER met2 ( -140 -2000 ) ( 140 2000 )
x[28], LAYER met2 ( -140 -2000 ) ( 140 2000 )
x[29], LAYER met2 ( -140 -2000 ) ( 140 2000 )
x[30], LAYER met3 ( -2000 -300 ) ( 2000 300 )
x[31], LAYER met2 ( -140 -2000 ) ( 140 2000 )
y, LAYER met3 ( -2000 -300 ) ( 2000 300 )
#S
p, LAYER met3 ( -2000 -300 ) ( 2000 300 )
#E
clk, LAYER met2 ( -140 -2000 ) ( 140 2000 )
rst, LAYER met2 ( -140 -2000 ) ( 140 2000 )

